class driver;

endclass;